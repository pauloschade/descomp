library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3;
			 opcodeSize: natural := 4
    );
   port (
          address : in std_logic_vector (addrWidth-1 DOWNTO 0);
          data : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;



architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  
tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(1) := STA & "000" & "000001000"; -- STA [0] @8

tmp(2) := LDI & "111" & "000000001"; -- LDI [7] $1

tmp(3) := STA & "111" & "000001001"; -- STA [7] @9

tmp(4) := LDI & "111" & "000001001"; -- LDI [7] $9

tmp(5) := STA & "111" & "000001110"; -- STA [7] @14

tmp(6) := STA & "111" & "000000010"; -- STA [7] @2

tmp(7) := STA & "111" & "000000011"; -- STA [7] @3

tmp(8) := STA & "111" & "000000100"; -- STA [7] @4

tmp(9) := STA & "111" & "000000101"; -- STA [7] @5

tmp(10) := STA & "111" & "000000110"; -- STA [7] @6

tmp(11) := STA & "111" & "000000111"; -- STA [7] @7

tmp(12) := STA & "000" & "111111111"; -- STA @511

tmp(13) := STA & "000" & "111111110"; -- STA @510

tmp(14) := LDA & "111" & "101100100"; -- LDA [7] @356

tmp(15) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(16) := JEQ & "000" & "001001000"; -- JEQ @72

tmp(17) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(18) := CEQ & "111" & "000001001"; -- CEQ [7] @9

tmp(19) := JEQ & "000" & "001010101"; -- JEQ @85

tmp(20) := LDA & "111" & "101100000"; -- LDA [7] @352

tmp(21) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(22) := JEQ & "000" & "000001110"; -- JEQ @14

tmp(23) := JSR & "000" & "010001010"; -- JSR @138

tmp(24) := LDA & "110" & "000001000"; -- LDA [6] @8

tmp(25) := STA & "110" & "100000001"; -- STA [6] @257

tmp(26) := JSR & "000" & "000011100"; -- JSR @28

tmp(27) := JMP & "000" & "000001110"; -- JMP @14

tmp(28) := STA & "000" & "111111111"; -- STA @511

tmp(29) := CEQ & "000" & "000001110"; -- CEQ [0] @14

tmp(30) := JEQ & "000" & "000100010"; -- JEQ @34

tmp(31) := SOMA & "000" & "000001001"; -- SOMA [0] @9

tmp(32) := STA & "000" & "100100000"; -- STA [0] @288

tmp(33) := RET & "000" & "000000000"; -- RET

tmp(34) := LDA & "000" & "000001000"; -- LDA [0] @8

tmp(35) := STA & "000" & "100100000"; -- STA [0] @288

tmp(36) := CEQ & "001" & "000001110"; -- CEQ [1] @14

tmp(37) := JEQ & "000" & "000101001"; -- JEQ @41

tmp(38) := SOMA & "001" & "000001001"; -- SOMA [1] @9

tmp(39) := STA & "001" & "100100001"; -- STA [1] @289

tmp(40) := RET & "000" & "000000000"; -- RET

tmp(41) := LDA & "001" & "000001000"; -- LDA [1] @8

tmp(42) := STA & "001" & "100100001"; -- STA [1] @289

tmp(43) := CEQ & "010" & "000001110"; -- CEQ [2] @14

tmp(44) := JEQ & "000" & "000110000"; -- JEQ @48

tmp(45) := SOMA & "010" & "000001001"; -- SOMA [2] @9

tmp(46) := STA & "010" & "100100010"; -- STA [2] @290

tmp(47) := RET & "000" & "000000000"; -- RET

tmp(48) := LDA & "010" & "000001000"; -- LDA [2] @8

tmp(49) := STA & "010" & "100100010"; -- STA [2] @290

tmp(50) := CEQ & "011" & "000001110"; -- CEQ [3] @14

tmp(51) := JEQ & "000" & "000110111"; -- JEQ @55

tmp(52) := SOMA & "011" & "000001001"; -- SOMA [3] @9

tmp(53) := STA & "011" & "100100011"; -- STA [3] @291

tmp(54) := RET & "000" & "000000000"; -- RET

tmp(55) := LDA & "011" & "000001000"; -- LDA [3] @8

tmp(56) := STA & "011" & "100100011"; -- STA [3] @291

tmp(57) := CEQ & "100" & "000001110"; -- CEQ [4] @14

tmp(58) := JEQ & "000" & "000111110"; -- JEQ @62

tmp(59) := SOMA & "100" & "000001001"; -- SOMA [4] @9

tmp(60) := STA & "100" & "100100100"; -- STA [4] @292

tmp(61) := RET & "000" & "000000000"; -- RET

tmp(62) := LDA & "100" & "000001000"; -- LDA [4] @8

tmp(63) := STA & "100" & "100100100"; -- STA [4] @292

tmp(64) := CEQ & "101" & "000001110"; -- CEQ [5] @14

tmp(65) := JEQ & "000" & "001000101"; -- JEQ @69

tmp(66) := SOMA & "101" & "000001001"; -- SOMA [5] @9

tmp(67) := STA & "101" & "100100101"; -- STA [5] @293

tmp(68) := RET & "000" & "000000000"; -- RET

tmp(69) := LDI & "110" & "000001001"; -- LDI [6] @9

tmp(70) := STA & "110" & "100000010"; -- STA [6] @258

tmp(71) := RET & "000" & "000000000"; -- RET

tmp(72) := LDI & "000" & "000000000"; -- LDI [0] $0

tmp(73) := LDI & "001" & "000000000"; -- LDI [1] $0

tmp(74) := LDI & "010" & "000000000"; -- LDI [2] $0

tmp(75) := LDI & "011" & "000000000"; -- LDI [3] $0

tmp(76) := LDI & "100" & "000000000"; -- LDI [4] $0

tmp(77) := LDI & "101" & "000000000"; -- LDI [5] $0

tmp(78) := STA & "000" & "100100000"; -- STA [0] @288

tmp(79) := STA & "001" & "100100001"; -- STA [1] @289

tmp(80) := STA & "010" & "100100010"; -- STA [2] @290

tmp(81) := STA & "011" & "100100011"; -- STA [3] @291

tmp(82) := STA & "100" & "100100100"; -- STA [4] @292

tmp(83) := STA & "101" & "100100101"; -- STA [5] @293

tmp(84) := JMP & "000" & "000001110"; -- JMP @14

tmp(85) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(86) := STA & "110" & "100100000"; -- STA [6] @288

tmp(87) := STA & "110" & "000000010"; -- STA [6] @2

tmp(88) := STA & "000" & "111111110"; -- STA @510

tmp(89) := LDI & "000" & "000000010"; -- LDI [0] $2

tmp(90) := STA & "000" & "100000000"; -- STA [0] @256

tmp(91) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(92) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(93) := JEQ & "000" & "001011011"; -- JEQ @91

tmp(94) := STA & "000" & "111111110"; -- STA @510

tmp(95) := LDI & "000" & "000000100"; -- LDI [0] $4

tmp(96) := STA & "000" & "100000000"; -- STA [0] @256

tmp(97) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(98) := STA & "110" & "100100001"; -- STA [6] @289

tmp(99) := STA & "110" & "000000011"; -- STA [6] @3

tmp(100) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(101) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(102) := JEQ & "000" & "001100100"; -- JEQ @100

tmp(103) := STA & "000" & "111111110"; -- STA @510

tmp(104) := LDI & "000" & "000001000"; -- LDI [0] $8

tmp(105) := STA & "000" & "100000000"; -- STA [0] @256

tmp(106) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(107) := STA & "110" & "100100010"; -- STA [6] @290

tmp(108) := STA & "110" & "000000100"; -- STA [6] @4

tmp(109) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(110) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(111) := JEQ & "000" & "001101101"; -- JEQ @109

tmp(112) := STA & "000" & "111111110"; -- STA @510

tmp(113) := LDI & "000" & "000010000"; -- LDI [0] $16

tmp(114) := STA & "000" & "100000000"; -- STA [0] @256

tmp(115) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(116) := STA & "110" & "100100011"; -- STA [6] @291

tmp(117) := STA & "110" & "000000101"; -- STA [6] @5

tmp(118) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(119) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(120) := JEQ & "000" & "001110110"; -- JEQ @118

tmp(121) := STA & "000" & "111111110"; -- STA @510

tmp(122) := LDI & "000" & "000100000"; -- LDI [0] $32

tmp(123) := STA & "000" & "100000000"; -- STA [0] @256

tmp(124) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(125) := STA & "110" & "100100100"; -- STA [6] @292

tmp(126) := STA & "110" & "000000110"; -- STA [6] @6

tmp(127) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(128) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(129) := JEQ & "000" & "001111111"; -- JEQ @127

tmp(130) := STA & "000" & "111111110"; -- STA @510

tmp(131) := LDI & "000" & "000000000"; -- LDI [0] $0

tmp(132) := STA & "000" & "100000000"; -- STA [0] @256

tmp(133) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(134) := STA & "110" & "100100101"; -- STA [6] @293

tmp(135) := STA & "110" & "000000111"; -- STA [6] @7

tmp(136) := STA & "000" & "111111110"; -- STA @510

tmp(137) := JMP & "000" & "001001000"; -- JMP @72

tmp(138) := STA & "000" & "111111111"; -- STA @511

tmp(139) := CEQ & "101" & "000000111"; -- CEQ [5] @7

tmp(140) := JEQ & "000" & "010001110"; -- JEQ @142

tmp(141) := RET & "000" & "000000000"; -- RET

tmp(142) := CEQ & "100" & "000000110"; -- CEQ [4] @6

tmp(143) := JEQ & "000" & "010010001"; -- JEQ @145

tmp(144) := RET & "000" & "000000000"; -- RET

tmp(145) := CEQ & "011" & "000000101"; -- CEQ [3] @5

tmp(146) := JEQ & "000" & "010010100"; -- JEQ @148

tmp(147) := RET & "000" & "000000000"; -- RET

tmp(148) := CEQ & "010" & "000000100"; -- CEQ [2] @4

tmp(149) := JEQ & "000" & "010010111"; -- JEQ @151

tmp(150) := RET & "000" & "000000000"; -- RET

tmp(151) := CEQ & "001" & "000000011"; -- CEQ [1] @3

tmp(152) := JEQ & "000" & "010011010"; -- JEQ @154

tmp(153) := RET & "000" & "000000000"; -- RET

tmp(154) := CEQ & "000" & "000000010"; -- CEQ [0] @2

tmp(155) := LDA & "110" & "000001001"; -- LDA [6] @9

tmp(156) := STA & "110" & "100000001"; -- STA [6] @257

tmp(157) := JEQ & "000" & "000001110"; -- JEQ @14

tmp(158) := RET & "000" & "000000000"; -- RET

  
--tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0
--
--tmp(1) := STA & "000" & "000001000"; -- STA [0] @8
--
--tmp(2) := LDI & "111" & "000000001"; -- LDI [7] $1
--
--tmp(3) := STA & "111" & "000001001"; -- STA [7] @9
--
--tmp(4) := LDI & "111" & "000001001"; -- LDI [7] $9
--
--tmp(5) := STA & "111" & "000001110"; -- STA [7] @14
--
--tmp(6) := STA & "000" & "111111111"; -- STA @511
--
--tmp(7) := STA & "000" & "111111110"; -- STA @510
--
--tmp(8) := LDA & "111" & "101100100"; -- LDA [7] @356
--
--tmp(9) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(10) := JEQ & "000" & "000111111"; -- JEQ @63
--
--tmp(11) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(12) := CEQ & "111" & "000001001"; -- CEQ [7] @9
--
--tmp(13) := JEQ & "000" & "001001100"; -- JEQ @76
--
--tmp(14) := LDA & "111" & "101100000"; -- LDA [7] @352
--
--tmp(15) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(16) := JEQ & "000" & "000001000"; -- JEQ @8
--
--tmp(17) := JSR & "000" & "000010011"; -- JSR @19
--
--tmp(18) := JMP & "000" & "000001000"; -- JMP @8
--
--tmp(19) := STA & "000" & "111111111"; -- STA @511
--
--tmp(20) := CEQ & "000" & "000001110"; -- CEQ [0] @14
--
--tmp(21) := JEQ & "000" & "000011001"; -- JEQ @25
--
--tmp(22) := SOMA & "000" & "000001001"; -- SOMA [0] @9
--
--tmp(23) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(24) := RET & "000" & "000000000"; -- RET
--
--tmp(25) := LDA & "000" & "000001000"; -- LDA [0] @8
--
--tmp(26) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(27) := CEQ & "001" & "000001110"; -- CEQ [1] @14
--
--tmp(28) := JEQ & "000" & "000100000"; -- JEQ @32
--
--tmp(29) := SOMA & "001" & "000001001"; -- SOMA [1] @9
--
--tmp(30) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(31) := RET & "000" & "000000000"; -- RET
--
--tmp(32) := LDA & "001" & "000001000"; -- LDA [1] @8
--
--tmp(33) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(34) := CEQ & "010" & "000001110"; -- CEQ [2] @14
--
--tmp(35) := JEQ & "000" & "000100111"; -- JEQ @39
--
--tmp(36) := SOMA & "010" & "000001001"; -- SOMA [2] @9
--
--tmp(37) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(38) := RET & "000" & "000000000"; -- RET
--
--tmp(39) := LDA & "010" & "000001000"; -- LDA [2] @8
--
--tmp(40) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(41) := CEQ & "011" & "000001110"; -- CEQ [3] @14
--
--tmp(42) := JEQ & "000" & "000101110"; -- JEQ @46
--
--tmp(43) := SOMA & "011" & "000001001"; -- SOMA [3] @9
--
--tmp(44) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(45) := RET & "000" & "000000000"; -- RET
--
--tmp(46) := LDA & "011" & "000001000"; -- LDA [3] @8
--
--tmp(47) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(48) := CEQ & "100" & "000001110"; -- CEQ [4] @14
--
--tmp(49) := JEQ & "000" & "000110101"; -- JEQ @53
--
--tmp(50) := SOMA & "100" & "000001001"; -- SOMA [4] @9
--
--tmp(51) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(52) := RET & "000" & "000000000"; -- RET
--
--tmp(53) := LDA & "100" & "000001000"; -- LDA [4] @8
--
--tmp(54) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(55) := CEQ & "101" & "000001110"; -- CEQ [5] @14
--
--tmp(56) := JEQ & "000" & "000111100"; -- JEQ @60
--
--tmp(57) := SOMA & "101" & "000001001"; -- SOMA [5] @9
--
--tmp(58) := STA & "101" & "100100101"; -- STA [5] @293
--
--tmp(59) := RET & "000" & "000000000"; -- RET
--
--tmp(60) := LDI & "110" & "000000001"; -- LDI [6] $1
--
--tmp(61) := STA & "110" & "100000010"; -- STA [6] @258
--
--tmp(62) := RET & "000" & "000000000"; -- RET
--
--tmp(63) := LDI & "000" & "000000000"; -- LDI [0] $0
--
--tmp(64) := LDI & "001" & "000000000"; -- LDI [1] $0
--
--tmp(65) := LDI & "010" & "000000000"; -- LDI [2] $0
--
--tmp(66) := LDI & "011" & "000000000"; -- LDI [3] $0
--
--tmp(67) := LDI & "100" & "000000000"; -- LDI [4] $0
--
--tmp(68) := LDI & "101" & "000000000"; -- LDI [5] $0
--
--tmp(69) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(70) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(71) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(72) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(73) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(74) := STA & "101" & "100100101"; -- STA [5] @293
--
--tmp(75) := JMP & "000" & "000001000"; -- JMP @8
--
--tmp(76) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(77) := STA & "110" & "100100000"; -- STA [6] @288
--
--tmp(78) := STA & "110" & "000000010"; -- STA [6] @2
--
--tmp(79) := STA & "000" & "111111110"; -- STA @510
--
--tmp(80) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(81) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(82) := JEQ & "000" & "001010000"; -- JEQ @80
--
--tmp(83) := STA & "000" & "111111110"; -- STA @510
--
--tmp(84) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(85) := STA & "110" & "100100001"; -- STA [6] @289
--
--tmp(86) := STA & "110" & "000000011"; -- STA [6] @3
--
--tmp(87) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(88) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(89) := JEQ & "000" & "001010111"; -- JEQ @87
--
--tmp(90) := STA & "000" & "111111110"; -- STA @510
--
--tmp(91) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(92) := STA & "110" & "100100010"; -- STA [6] @290
--
--tmp(93) := STA & "110" & "000000100"; -- STA [6] @4
--
--tmp(94) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(95) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(96) := JEQ & "000" & "001011110"; -- JEQ @94
--
--tmp(97) := STA & "000" & "111111110"; -- STA @510
--
--tmp(98) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(99) := STA & "110" & "100100011"; -- STA [6] @291
--
--tmp(100) := STA & "110" & "000000101"; -- STA [6] @5
--
--tmp(101) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(102) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(103) := JEQ & "000" & "001100101"; -- JEQ @101
--
--tmp(104) := STA & "000" & "111111110"; -- STA @510
--
--tmp(105) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(106) := STA & "110" & "100100100"; -- STA [6] @292
--
--tmp(107) := STA & "110" & "000000110"; -- STA [6] @6
--
--tmp(108) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(109) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(110) := JEQ & "000" & "001101100"; -- JEQ @108
--
--tmp(111) := STA & "000" & "111111110"; -- STA @510
--
--tmp(112) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(113) := STA & "110" & "100100101"; -- STA [6] @293
--
--tmp(114) := STA & "110" & "000000111"; -- STA [6] @7
--
--tmp(115) := STA & "000" & "111111110"; -- STA @510
--
--tmp(116) := JMP & "000" & "000111111"; -- JMP @63



        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    data <= memROM (to_integer(unsigned(address)));
end architecture;