library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3;
			 opcodeSize: natural := 4
    );
   port (
          address : in std_logic_vector (addrWidth-1 DOWNTO 0);
          data : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;



architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDB  : std_logic_vector(3 downto 0) := "1011";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
<<<<<<< Updated upstream
			
tmp(0) := LDI & "111" & "000000000"; -- LDI R7 $0
=======
  
tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0
>>>>>>> Stashed changes

tmp(1) := STA & "000" & "000001000"; -- STA R0 @MEM0

tmp(2) := LDI & "111" & "000000001"; -- LDI R7 $1

tmp(3) := STA & "111" & "000001001"; -- STA R7 @MEM1

tmp(4) := LDI & "111" & "000001001"; -- LDI R7 $9

<<<<<<< Updated upstream
tmp(5) := STA & "111" & "000001110"; -- STA R7 @MEM9
=======
tmp(5) := STA & "111" & "000010000"; -- STA [7] @16
>>>>>>> Stashed changes

tmp(6) := LDI & "000" & "000000000"; -- LDI R0 $0

tmp(7) := LDI & "001" & "000000000"; -- LDI R1 $0

tmp(8) := LDI & "010" & "000000000"; -- LDI R2 $0

tmp(9) := LDI & "011" & "000000000"; -- LDI R3 $0

tmp(10) := LDI & "100" & "000000000"; -- LDI R4 $0

tmp(11) := LDA & "111" & "101100000"; -- LDA R7 @KEY0

<<<<<<< Updated upstream
tmp(12) := CEQ & "111" & "000000000"; -- CEQ R7 @0

tmp(13) := JEQ & "000" & "000001011"; -- JEQ @11

tmp(14) := JSR & "000" & "000010000"; -- JSR @16

tmp(15) := JMP & "000" & "000001011"; -- JMP @11

tmp(16) := STA & "000" & "111111111"; -- STA @clr_KEY0

tmp(17) := CEQ & "000" & "000001110"; -- CEQ R0 @MEM9

tmp(18) := JEQ & "000" & "000010110"; -- JEQ @22

tmp(19) := SOMA & "000" & "000001001"; -- SOMA R0 @MEM1

tmp(20) := STA & "000" & "100100000"; -- STA R0 @HEX0

tmp(21) := RET & "000" & "000000000"; -- RET

tmp(22) := LDA & "000" & "000001000"; -- LDA R0 $MEM0

tmp(23) := STA & "000" & "100100000"; -- STA R0 @HEX0

tmp(24) := CEQ & "001" & "000001110"; -- CEQ R1 @MEM9

tmp(25) := JEQ & "000" & "000011101"; -- JEQ @29

tmp(26) := SOMA & "001" & "000001001"; -- SOMA R1 @MEM1

tmp(27) := STA & "001" & "100100001"; -- STA R1 @HEX1

tmp(28) := RET & "000" & "000000000"; -- RET

tmp(29) := LDA & "001" & "000001000"; -- LDA R1 $MEM0

tmp(30) := STA & "001" & "100100001"; -- STA R1 @HEX1

tmp(31) := CEQ & "010" & "000001110"; -- CEQ R2 @MEM9

tmp(32) := JEQ & "000" & "000100100"; -- JEQ @36

tmp(33) := SOMA & "010" & "000001001"; -- SOMA R2 @MEM1

tmp(34) := STA & "010" & "100100010"; -- STA R2 @HEX2

tmp(35) := RET & "000" & "000000000"; -- RET

tmp(36) := LDA & "010" & "000001000"; -- LDA R2 $MEM0

tmp(37) := STA & "010" & "100100010"; -- STA R2 @HEX2

tmp(38) := CEQ & "011" & "000001110"; -- CEQ R3 @MEM9

tmp(39) := JEQ & "000" & "000100100"; -- JEQ @36

tmp(40) := SOMA & "011" & "000001001"; -- SOMA R3 @MEM1

tmp(41) := STA & "011" & "100100011"; -- STA R3 @HEX3
=======
tmp(12) := LDI & "111" & "010000000"; -- LDI [7] $128

tmp(13) := STA & "111" & "000001100"; -- STA [7] @12

tmp(14) := STA & "000" & "111111111"; -- STA @511

tmp(15) := STA & "000" & "111111110"; -- STA @510

tmp(16) := JMP & "000" & "001001011"; -- JMP @75

tmp(17) := LDA & "111" & "101100100"; -- LDA [7] @356

tmp(18) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(19) := JEQ & "000" & "001001011"; -- JEQ @75

tmp(20) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(21) := CEQ & "111" & "000001001"; -- CEQ [7] @9

tmp(22) := JEQ & "000" & "001100010"; -- JEQ @98

tmp(23) := LDA & "111" & "101100000"; -- LDA [7] @352

tmp(24) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(25) := JEQ & "000" & "000010001"; -- JEQ @17

tmp(26) := JSR & "000" & "010101000"; -- JSR @168

tmp(27) := LDA & "110" & "000001000"; -- LDA [6] @8

tmp(28) := STA & "110" & "100000001"; -- STA [6] @257

tmp(29) := JSR & "000" & "000011111"; -- JSR @31

tmp(30) := JMP & "000" & "000010001"; -- JMP @17

tmp(31) := STA & "000" & "111111111"; -- STA @511

tmp(32) := CEQ & "000" & "000010000"; -- CEQ [0] @16

tmp(33) := JEQ & "000" & "000100101"; -- JEQ @37

tmp(34) := SOMA & "000" & "000001001"; -- SOMA [0] @9

tmp(35) := STA & "000" & "100100000"; -- STA [0] @288

tmp(36) := RET & "000" & "000000000"; -- RET

tmp(37) := LDA & "000" & "000001000"; -- LDA [0] @8

tmp(38) := STA & "000" & "100100000"; -- STA [0] @288

tmp(39) := CEQ & "001" & "000010000"; -- CEQ [1] @16

tmp(40) := JEQ & "000" & "000101100"; -- JEQ @44

tmp(41) := SOMA & "001" & "000001001"; -- SOMA [1] @9

tmp(42) := STA & "001" & "100100001"; -- STA [1] @289

tmp(43) := RET & "000" & "000000000"; -- RET

tmp(44) := LDA & "001" & "000001000"; -- LDA [1] @8

tmp(45) := STA & "001" & "100100001"; -- STA [1] @289

tmp(46) := CEQ & "010" & "000010000"; -- CEQ [2] @16

tmp(47) := JEQ & "000" & "000110011"; -- JEQ @51

tmp(48) := SOMA & "010" & "000001001"; -- SOMA [2] @9

tmp(49) := STA & "010" & "100100010"; -- STA [2] @290

tmp(50) := RET & "000" & "000000000"; -- RET

tmp(51) := LDA & "010" & "000001000"; -- LDA [2] @8

tmp(52) := STA & "010" & "100100010"; -- STA [2] @290

tmp(53) := CEQ & "011" & "000010000"; -- CEQ [3] @16

tmp(54) := JEQ & "000" & "000111010"; -- JEQ @58

tmp(55) := SOMA & "011" & "000001001"; -- SOMA [3] @9

tmp(56) := STA & "011" & "100100011"; -- STA [3] @291

tmp(57) := RET & "000" & "000000000"; -- RET

tmp(58) := LDA & "011" & "000001000"; -- LDA [3] @8

tmp(59) := STA & "011" & "100100011"; -- STA [3] @291

tmp(60) := CEQ & "100" & "000010000"; -- CEQ [4] @16

tmp(61) := JEQ & "000" & "001000001"; -- JEQ @65

tmp(62) := SOMA & "100" & "000001001"; -- SOMA [4] @9

tmp(63) := STA & "100" & "100100100"; -- STA [4] @292

tmp(64) := RET & "000" & "000000000"; -- RET

tmp(65) := LDA & "100" & "000001000"; -- LDA [4] @8

tmp(66) := STA & "100" & "100100100"; -- STA [4] @292

tmp(67) := CEQ & "101" & "000010000"; -- CEQ [5] @16

tmp(68) := JEQ & "000" & "001001000"; -- JEQ @72

tmp(69) := SOMA & "101" & "000001001"; -- SOMA [5] @9

tmp(70) := STA & "101" & "100100101"; -- STA [5] @293

tmp(71) := RET & "000" & "000000000"; -- RET

tmp(72) := LDI & "110" & "000001001"; -- LDI [6] @9

tmp(73) := STA & "110" & "100000010"; -- STA [6] @258

tmp(74) := RET & "000" & "000000000"; -- RET

tmp(75) := LDI & "000" & "000000000"; -- LDI [0] $0

tmp(76) := LDI & "001" & "000000000"; -- LDI [1] $0

tmp(77) := LDI & "010" & "000000000"; -- LDI [2] $0

tmp(78) := LDI & "011" & "000000000"; -- LDI [3] $0

tmp(79) := LDI & "100" & "000000000"; -- LDI [4] $0

tmp(80) := LDI & "101" & "000000000"; -- LDI [5] $0

tmp(81) := JSR & "000" & "001010011"; -- JSR @83

tmp(82) := JMP & "000" & "000010001"; -- JMP @17

tmp(83) := STA & "000" & "100100000"; -- STA [0] @288

tmp(84) := STA & "001" & "100100001"; -- STA [1] @289

tmp(85) := STA & "010" & "100100010"; -- STA [2] @290

tmp(86) := STA & "011" & "100100011"; -- STA [3] @291

tmp(87) := STA & "100" & "100100100"; -- STA [4] @292

tmp(88) := STA & "101" & "100100101"; -- STA [5] @293

tmp(89) := RET & "000" & "000000000"; -- RET

tmp(90) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(91) := STA & "111" & "100100000"; -- STA [7] @288

tmp(92) := STA & "111" & "100100001"; -- STA [7] @289

tmp(93) := STA & "111" & "100100010"; -- STA [7] @290

tmp(94) := STA & "111" & "100100011"; -- STA [7] @291

tmp(95) := STA & "111" & "100100100"; -- STA [7] @292

tmp(96) := STA & "111" & "100100101"; -- STA [7] @293

tmp(97) := RET & "000" & "000000000"; -- RET

tmp(98) := JSR & "000" & "001011010"; -- JSR @90

tmp(99) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(100) := LDA & "111" & "000010000"; -- LDA [7] @16

tmp(101) := JSR & "000" & "010111100"; -- JSR @188

tmp(102) := STA & "110" & "100100000"; -- STA [6] @288

tmp(103) := STA & "110" & "000000010"; -- STA [6] @2

tmp(104) := STA & "000" & "111111110"; -- STA @510

tmp(105) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(106) := STA & "111" & "100000000"; -- STA [7] @256

tmp(107) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(108) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(109) := JEQ & "000" & "001101011"; -- JEQ @107

tmp(110) := STA & "000" & "111111110"; -- STA @510

tmp(111) := LDI & "111" & "000000100"; -- LDI [7] $4

tmp(112) := STA & "111" & "100000000"; -- STA [7] @256

tmp(113) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(114) := LDA & "111" & "000010000"; -- LDA [7] @16

tmp(115) := JSR & "000" & "010111100"; -- JSR @188

tmp(116) := STA & "110" & "100100001"; -- STA [6] @289

tmp(117) := STA & "110" & "000000011"; -- STA [6] @3

tmp(118) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(119) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(120) := JEQ & "000" & "001110110"; -- JEQ @118

tmp(121) := STA & "000" & "111111110"; -- STA @510

tmp(122) := LDI & "111" & "000001000"; -- LDI [7] $8

tmp(123) := STA & "111" & "100000000"; -- STA [7] @256

tmp(124) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(125) := LDA & "111" & "000010000"; -- LDA [7] @16

tmp(126) := JSR & "000" & "010111100"; -- JSR @188

tmp(127) := STA & "110" & "100100010"; -- STA [6] @290

tmp(128) := STA & "110" & "000000100"; -- STA [6] @4

tmp(129) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(130) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(131) := JEQ & "000" & "010000001"; -- JEQ @129

tmp(132) := STA & "000" & "111111110"; -- STA @510

tmp(133) := LDI & "111" & "000010000"; -- LDI [7] $16

tmp(134) := STA & "111" & "100000000"; -- STA [7] @256

tmp(135) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(136) := LDA & "111" & "000010000"; -- LDA [7] @16

tmp(137) := JSR & "000" & "010111100"; -- JSR @188

tmp(138) := STA & "110" & "100100011"; -- STA [6] @291

tmp(139) := STA & "110" & "000000101"; -- STA [6] @5

tmp(140) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(141) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(142) := JEQ & "000" & "010001100"; -- JEQ @140

tmp(143) := STA & "000" & "111111110"; -- STA @510

tmp(144) := LDI & "111" & "000100000"; -- LDI [7] $32

tmp(145) := STA & "111" & "100000000"; -- STA [7] @256

tmp(146) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(147) := LDA & "111" & "000010000"; -- LDA [7] @16

tmp(148) := JSR & "000" & "010111100"; -- JSR @188

tmp(149) := STA & "110" & "100100100"; -- STA [6] @292

tmp(150) := STA & "110" & "000000110"; -- STA [6] @6

tmp(151) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(152) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(153) := JEQ & "000" & "010010111"; -- JEQ @151

tmp(154) := STA & "000" & "111111110"; -- STA @510

tmp(155) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(156) := STA & "111" & "100000000"; -- STA [7] @256

tmp(157) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(158) := LDA & "111" & "000010000"; -- LDA [7] @16

tmp(159) := JSR & "000" & "010111100"; -- JSR @188

tmp(160) := STA & "110" & "100100101"; -- STA [6] @293

tmp(161) := STA & "110" & "000000111"; -- STA [6] @7

tmp(162) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(163) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(164) := JEQ & "000" & "010100010"; -- JEQ @162

tmp(165) := STA & "000" & "111111110"; -- STA @510

tmp(166) := JSR & "000" & "001010011"; -- JSR @83

tmp(167) := JMP & "000" & "000010001"; -- JMP @17

tmp(168) := CEQ & "101" & "000000111"; -- CEQ [5] @7

tmp(169) := JEQ & "000" & "010101011"; -- JEQ @171

tmp(170) := RET & "000" & "000000000"; -- RET

tmp(171) := CEQ & "100" & "000000110"; -- CEQ [4] @6

tmp(172) := JEQ & "000" & "010101110"; -- JEQ @174

tmp(173) := RET & "000" & "000000000"; -- RET

tmp(174) := CEQ & "011" & "000000101"; -- CEQ [3] @5

tmp(175) := JEQ & "000" & "010110001"; -- JEQ @177

tmp(176) := RET & "000" & "000000000"; -- RET

tmp(177) := CEQ & "010" & "000000100"; -- CEQ [2] @4

tmp(178) := JEQ & "000" & "010110100"; -- JEQ @180

tmp(179) := RET & "000" & "000000000"; -- RET

tmp(180) := CEQ & "001" & "000000011"; -- CEQ [1] @3

tmp(181) := JEQ & "000" & "010110111"; -- JEQ @183

tmp(182) := RET & "000" & "000000000"; -- RET

tmp(183) := CEQ & "000" & "000000010"; -- CEQ [0] @2

tmp(184) := LDA & "110" & "000001001"; -- LDA [6] @9

tmp(185) := STA & "110" & "100000001"; -- STA [6] @257

tmp(186) := JEQ & "000" & "000010001"; -- JEQ @17

tmp(187) := RET & "000" & "000000000"; -- RET

tmp(188) := STA & "110" & "000001101"; -- STA [6] @13

tmp(189) := STA & "111" & "000001110"; -- STA [7] @14

tmp(190) := SUB & "111" & "000001101"; -- SUB [7] @13

tmp(191) := ANDB & "111" & "000001100"; -- ANDB [7] @12

tmp(192) := CEQ & "111" & "000001100"; -- CEQ [7] @12

tmp(193) := JEQ & "000" & "011000100"; -- JEQ @196

tmp(194) := STA & "111" & "000001000"; -- STA [7] @8

tmp(195) := RET & "000" & "000000000"; -- RET

tmp(196) := STA & "111" & "000001001"; -- STA [7] @9

tmp(197) := LDA & "110" & "000001110"; -- LDA [6] @14

tmp(198) := RET & "000" & "000000000"; -- RET

  
--tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0
--
--tmp(1) := STA & "000" & "000001000"; -- STA [0] @8
--
--tmp(2) := LDI & "111" & "000000001"; -- LDI [7] $1
--
--tmp(3) := STA & "111" & "000001001"; -- STA [7] @9
--
--tmp(4) := LDI & "111" & "000001001"; -- LDI [7] $9
--
--tmp(5) := STA & "111" & "000001110"; -- STA [7] @14
--
--tmp(6) := STA & "000" & "111111111"; -- STA @511
--
--tmp(7) := STA & "000" & "111111110"; -- STA @510
--
--tmp(8) := LDA & "111" & "101100100"; -- LDA [7] @356
--
--tmp(9) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(10) := JEQ & "000" & "000111111"; -- JEQ @63
--
--tmp(11) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(12) := CEQ & "111" & "000001001"; -- CEQ [7] @9
--
--tmp(13) := JEQ & "000" & "001001100"; -- JEQ @76
--
--tmp(14) := LDA & "111" & "101100000"; -- LDA [7] @352
--
--tmp(15) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(16) := JEQ & "000" & "000001000"; -- JEQ @8
--
--tmp(17) := JSR & "000" & "000010011"; -- JSR @19
--
--tmp(18) := JMP & "000" & "000001000"; -- JMP @8
--
--tmp(19) := STA & "000" & "111111111"; -- STA @511
--
--tmp(20) := CEQ & "000" & "000001110"; -- CEQ [0] @14
--
--tmp(21) := JEQ & "000" & "000011001"; -- JEQ @25
--
--tmp(22) := SOMA & "000" & "000001001"; -- SOMA [0] @9
--
--tmp(23) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(24) := RET & "000" & "000000000"; -- RET
--
--tmp(25) := LDA & "000" & "000001000"; -- LDA [0] @8
--
--tmp(26) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(27) := CEQ & "001" & "000001110"; -- CEQ [1] @14
--
--tmp(28) := JEQ & "000" & "000100000"; -- JEQ @32
--
--tmp(29) := SOMA & "001" & "000001001"; -- SOMA [1] @9
--
--tmp(30) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(31) := RET & "000" & "000000000"; -- RET
--
--tmp(32) := LDA & "001" & "000001000"; -- LDA [1] @8
--
--tmp(33) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(34) := CEQ & "010" & "000001110"; -- CEQ [2] @14
--
--tmp(35) := JEQ & "000" & "000100111"; -- JEQ @39
--
--tmp(36) := SOMA & "010" & "000001001"; -- SOMA [2] @9
--
--tmp(37) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(38) := RET & "000" & "000000000"; -- RET
--
--tmp(39) := LDA & "010" & "000001000"; -- LDA [2] @8
--
--tmp(40) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(41) := CEQ & "011" & "000001110"; -- CEQ [3] @14
--
--tmp(42) := JEQ & "000" & "000101110"; -- JEQ @46
--
--tmp(43) := SOMA & "011" & "000001001"; -- SOMA [3] @9
--
--tmp(44) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(45) := RET & "000" & "000000000"; -- RET
--
--tmp(46) := LDA & "011" & "000001000"; -- LDA [3] @8
--
--tmp(47) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(48) := CEQ & "100" & "000001110"; -- CEQ [4] @14
--
--tmp(49) := JEQ & "000" & "000110101"; -- JEQ @53
--
--tmp(50) := SOMA & "100" & "000001001"; -- SOMA [4] @9
--
--tmp(51) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(52) := RET & "000" & "000000000"; -- RET
--
--tmp(53) := LDA & "100" & "000001000"; -- LDA [4] @8
--
--tmp(54) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(55) := CEQ & "101" & "000001110"; -- CEQ [5] @14
--
--tmp(56) := JEQ & "000" & "000111100"; -- JEQ @60
--
--tmp(57) := SOMA & "101" & "000001001"; -- SOMA [5] @9
--
--tmp(58) := STA & "101" & "100100101"; -- STA [5] @293
--
--tmp(59) := RET & "000" & "000000000"; -- RET
--
--tmp(60) := LDI & "110" & "000000001"; -- LDI [6] $1
--
--tmp(61) := STA & "110" & "100000010"; -- STA [6] @258
--
--tmp(62) := RET & "000" & "000000000"; -- RET
--
--tmp(63) := LDI & "000" & "000000000"; -- LDI [0] $0
--
--tmp(64) := LDI & "001" & "000000000"; -- LDI [1] $0
--
--tmp(65) := LDI & "010" & "000000000"; -- LDI [2] $0
--
--tmp(66) := LDI & "011" & "000000000"; -- LDI [3] $0
--
--tmp(67) := LDI & "100" & "000000000"; -- LDI [4] $0
--
--tmp(68) := LDI & "101" & "000000000"; -- LDI [5] $0
--
--tmp(69) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(70) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(71) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(72) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(73) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(74) := STA & "101" & "100100101"; -- STA [5] @293
--
--tmp(75) := JMP & "000" & "000001000"; -- JMP @8
--
--tmp(76) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(77) := STA & "110" & "100100000"; -- STA [6] @288
--
--tmp(78) := STA & "110" & "000000010"; -- STA [6] @2
--
--tmp(79) := STA & "000" & "111111110"; -- STA @510
--
--tmp(80) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(81) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(82) := JEQ & "000" & "001010000"; -- JEQ @80
--
--tmp(83) := STA & "000" & "111111110"; -- STA @510
--
--tmp(84) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(85) := STA & "110" & "100100001"; -- STA [6] @289
--
--tmp(86) := STA & "110" & "000000011"; -- STA [6] @3
--
--tmp(87) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(88) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(89) := JEQ & "000" & "001010111"; -- JEQ @87
--
--tmp(90) := STA & "000" & "111111110"; -- STA @510
--
--tmp(91) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(92) := STA & "110" & "100100010"; -- STA [6] @290
--
--tmp(93) := STA & "110" & "000000100"; -- STA [6] @4
--
--tmp(94) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(95) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(96) := JEQ & "000" & "001011110"; -- JEQ @94
--
--tmp(97) := STA & "000" & "111111110"; -- STA @510
--
--tmp(98) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(99) := STA & "110" & "100100011"; -- STA [6] @291
--
--tmp(100) := STA & "110" & "000000101"; -- STA [6] @5
--
--tmp(101) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(102) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(103) := JEQ & "000" & "001100101"; -- JEQ @101
--
--tmp(104) := STA & "000" & "111111110"; -- STA @510
--
--tmp(105) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(106) := STA & "110" & "100100100"; -- STA [6] @292
--
--tmp(107) := STA & "110" & "000000110"; -- STA [6] @6
--
--tmp(108) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(109) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(110) := JEQ & "000" & "001101100"; -- JEQ @108
--
--tmp(111) := STA & "000" & "111111110"; -- STA @510
--
--tmp(112) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(113) := STA & "110" & "100100101"; -- STA [6] @293
--
--tmp(114) := STA & "110" & "000000111"; -- STA [6] @7
--
--tmp(115) := STA & "000" & "111111110"; -- STA @510
--
--tmp(116) := JMP & "000" & "000111111"; -- JMP @63
>>>>>>> Stashed changes

tmp(42) := RET & "000" & "000000000"; -- RET


		  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    data <= memROM (to_integer(unsigned(address)));
end architecture;