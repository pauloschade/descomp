library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3;
			 opcodeSize: natural := 4
    );
   port (
          address : in std_logic_vector (addrWidth-1 DOWNTO 0);
          data : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;



architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
  

tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(1) := STA & "000" & "000001000"; -- STA [0] @8

tmp(2) := LDI & "111" & "000000001"; -- LDI [7] $1

tmp(3) := STA & "111" & "000001001"; -- STA [7] @9

tmp(4) := LDI & "111" & "000001001"; -- LDI [7] $9

tmp(5) := STA & "111" & "000001110"; -- STA [7] @14

tmp(6) := STA & "000" & "111111111"; -- STA @511

tmp(7) := STA & "000" & "111111110"; -- STA @510

tmp(8) := LDA & "111" & "101100100"; -- LDA [7] @356

tmp(9) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(10) := JEQ & "000" & "001000000"; -- JEQ @64

tmp(11) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(12) := CEQ & "111" & "000001001"; -- CEQ [7] @9

tmp(13) := JEQ & "000" & "001001101"; -- JEQ @77

tmp(14) := LDA & "111" & "101100000"; -- LDA [7] @352

tmp(15) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(16) := JEQ & "000" & "000001000"; -- JEQ @8

tmp(17) := JSR & "000" & "001110110"; -- JSR @118

tmp(18) := JSR & "000" & "000010100"; -- JSR @20

tmp(19) := JMP & "000" & "000001000"; -- JMP @8

tmp(20) := STA & "000" & "111111111"; -- STA @511

tmp(21) := CEQ & "000" & "000001110"; -- CEQ [0] @14

tmp(22) := JEQ & "000" & "000011010"; -- JEQ @26

tmp(23) := SOMA & "000" & "000001001"; -- SOMA [0] @9

tmp(24) := STA & "000" & "100100000"; -- STA [0] @288

tmp(25) := RET & "000" & "000000000"; -- RET

tmp(26) := LDA & "000" & "000001000"; -- LDA [0] @8

tmp(27) := STA & "000" & "100100000"; -- STA [0] @288

tmp(28) := CEQ & "001" & "000001110"; -- CEQ [1] @14

tmp(29) := JEQ & "000" & "000100001"; -- JEQ @33

tmp(30) := SOMA & "001" & "000001001"; -- SOMA [1] @9

tmp(31) := STA & "001" & "100100001"; -- STA [1] @289

tmp(32) := RET & "000" & "000000000"; -- RET

tmp(33) := LDA & "001" & "000001000"; -- LDA [1] @8

tmp(34) := STA & "001" & "100100001"; -- STA [1] @289

tmp(35) := CEQ & "010" & "000001110"; -- CEQ [2] @14

tmp(36) := JEQ & "000" & "000101000"; -- JEQ @40

tmp(37) := SOMA & "010" & "000001001"; -- SOMA [2] @9

tmp(38) := STA & "010" & "100100010"; -- STA [2] @290

tmp(39) := RET & "000" & "000000000"; -- RET

tmp(40) := LDA & "010" & "000001000"; -- LDA [2] @8

tmp(41) := STA & "010" & "100100010"; -- STA [2] @290

tmp(42) := CEQ & "011" & "000001110"; -- CEQ [3] @14

tmp(43) := JEQ & "000" & "000101111"; -- JEQ @47

tmp(44) := SOMA & "011" & "000001001"; -- SOMA [3] @9

tmp(45) := STA & "011" & "100100011"; -- STA [3] @291

tmp(46) := RET & "000" & "000000000"; -- RET

tmp(47) := LDA & "011" & "000001000"; -- LDA [3] @8

tmp(48) := STA & "011" & "100100011"; -- STA [3] @291

tmp(49) := CEQ & "100" & "000001110"; -- CEQ [4] @14

tmp(50) := JEQ & "000" & "000110110"; -- JEQ @54

tmp(51) := SOMA & "100" & "000001001"; -- SOMA [4] @9

tmp(52) := STA & "100" & "100100100"; -- STA [4] @292

tmp(53) := RET & "000" & "000000000"; -- RET

tmp(54) := LDA & "100" & "000001000"; -- LDA [4] @8

tmp(55) := STA & "100" & "100100100"; -- STA [4] @292

tmp(56) := CEQ & "101" & "000001110"; -- CEQ [5] @14

tmp(57) := JEQ & "000" & "000111101"; -- JEQ @61

tmp(58) := SOMA & "101" & "000001001"; -- SOMA [5] @9

tmp(59) := STA & "101" & "100100101"; -- STA [5] @293

tmp(60) := RET & "000" & "000000000"; -- RET

tmp(61) := LDI & "110" & "000000001"; -- LDI [6] $1

tmp(62) := STA & "110" & "100000010"; -- STA [6] @258

tmp(63) := RET & "000" & "000000000"; -- RET

tmp(64) := LDI & "000" & "000000000"; -- LDI [0] $0

tmp(65) := LDI & "001" & "000000000"; -- LDI [1] $0

tmp(66) := LDI & "010" & "000000000"; -- LDI [2] $0

tmp(67) := LDI & "011" & "000000000"; -- LDI [3] $0

tmp(68) := LDI & "100" & "000000000"; -- LDI [4] $0

tmp(69) := LDI & "101" & "000000000"; -- LDI [5] $0

tmp(70) := STA & "000" & "100100000"; -- STA [0] @288

tmp(71) := STA & "001" & "100100001"; -- STA [1] @289

tmp(72) := STA & "010" & "100100010"; -- STA [2] @290

tmp(73) := STA & "011" & "100100011"; -- STA [3] @291

tmp(74) := STA & "100" & "100100100"; -- STA [4] @292

tmp(75) := STA & "101" & "100100101"; -- STA [5] @293

tmp(76) := JMP & "000" & "000001000"; -- JMP @8

tmp(77) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(78) := STA & "110" & "100100000"; -- STA [6] @288

tmp(79) := STA & "110" & "000000010"; -- STA [6] @2

tmp(80) := STA & "000" & "111111110"; -- STA @510

tmp(81) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(82) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(83) := JEQ & "000" & "001010001"; -- JEQ @81

tmp(84) := STA & "000" & "111111110"; -- STA @510

tmp(85) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(86) := STA & "110" & "100100001"; -- STA [6] @289

tmp(87) := STA & "110" & "000000011"; -- STA [6] @3

tmp(88) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(89) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(90) := JEQ & "000" & "001011000"; -- JEQ @88

tmp(91) := STA & "000" & "111111110"; -- STA @510

tmp(92) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(93) := STA & "110" & "100100010"; -- STA [6] @290

tmp(94) := STA & "110" & "000000100"; -- STA [6] @4

tmp(95) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(96) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(97) := JEQ & "000" & "001011111"; -- JEQ @95

tmp(98) := STA & "000" & "111111110"; -- STA @510

tmp(99) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(100) := STA & "110" & "100100011"; -- STA [6] @291

tmp(101) := STA & "110" & "000000101"; -- STA [6] @5

tmp(102) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(103) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(104) := JEQ & "000" & "001100110"; -- JEQ @102

tmp(105) := STA & "000" & "111111110"; -- STA @510

tmp(106) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(107) := STA & "110" & "100100100"; -- STA [6] @292

tmp(108) := STA & "110" & "000000110"; -- STA [6] @6

tmp(109) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(110) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(111) := JEQ & "000" & "001101101"; -- JEQ @109

tmp(112) := STA & "000" & "111111110"; -- STA @510

tmp(113) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(114) := STA & "110" & "100100101"; -- STA [6] @293

tmp(115) := STA & "110" & "000000111"; -- STA [6] @7

tmp(116) := STA & "000" & "111111110"; -- STA @510

tmp(117) := JMP & "000" & "001000000"; -- JMP @64

tmp(118) := STA & "000" & "111111111"; -- STA @511

tmp(119) := CEQ & "101" & "000000111"; -- CEQ [5] @7

tmp(120) := JEQ & "000" & "001111010"; -- JEQ @122

tmp(121) := RET & "000" & "000000000"; -- RET

tmp(122) := CEQ & "100" & "000000110"; -- CEQ [4] @6

tmp(123) := JEQ & "000" & "001111101"; -- JEQ @125

tmp(124) := RET & "000" & "000000000"; -- RET

tmp(125) := CEQ & "011" & "000000101"; -- CEQ [3] @5

tmp(126) := JEQ & "000" & "010000000"; -- JEQ @128

tmp(127) := RET & "000" & "000000000"; -- RET

tmp(128) := CEQ & "010" & "000000100"; -- CEQ [2] @4

tmp(129) := JEQ & "000" & "010000011"; -- JEQ @131

tmp(130) := RET & "000" & "000000000"; -- RET

tmp(131) := CEQ & "001" & "000000011"; -- CEQ [1] @3

tmp(132) := JEQ & "000" & "010000110"; -- JEQ @134

tmp(133) := RET & "000" & "000000000"; -- RET

tmp(134) := CEQ & "000" & "000000010"; -- CEQ [0] @2

tmp(135) := JEQ & "000" & "000001000"; -- JEQ @8

tmp(136) := RET & "000" & "000000000"; -- RET


  
--tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0
--
--tmp(1) := STA & "000" & "000001000"; -- STA [0] @8
--
--tmp(2) := LDI & "111" & "000000001"; -- LDI [7] $1
--
--tmp(3) := STA & "111" & "000001001"; -- STA [7] @9
--
--tmp(4) := LDI & "111" & "000001001"; -- LDI [7] $9
--
--tmp(5) := STA & "111" & "000001110"; -- STA [7] @14
--
--tmp(6) := STA & "000" & "111111111"; -- STA @511
--
--tmp(7) := STA & "000" & "111111110"; -- STA @510
--
--tmp(8) := LDA & "111" & "101100100"; -- LDA [7] @356
--
--tmp(9) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(10) := JEQ & "000" & "000111111"; -- JEQ @63
--
--tmp(11) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(12) := CEQ & "111" & "000001001"; -- CEQ [7] @9
--
--tmp(13) := JEQ & "000" & "001001100"; -- JEQ @76
--
--tmp(14) := LDA & "111" & "101100000"; -- LDA [7] @352
--
--tmp(15) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(16) := JEQ & "000" & "000001000"; -- JEQ @8
--
--tmp(17) := JSR & "000" & "000010011"; -- JSR @19
--
--tmp(18) := JMP & "000" & "000001000"; -- JMP @8
--
--tmp(19) := STA & "000" & "111111111"; -- STA @511
--
--tmp(20) := CEQ & "000" & "000001110"; -- CEQ [0] @14
--
--tmp(21) := JEQ & "000" & "000011001"; -- JEQ @25
--
--tmp(22) := SOMA & "000" & "000001001"; -- SOMA [0] @9
--
--tmp(23) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(24) := RET & "000" & "000000000"; -- RET
--
--tmp(25) := LDA & "000" & "000001000"; -- LDA [0] @8
--
--tmp(26) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(27) := CEQ & "001" & "000001110"; -- CEQ [1] @14
--
--tmp(28) := JEQ & "000" & "000100000"; -- JEQ @32
--
--tmp(29) := SOMA & "001" & "000001001"; -- SOMA [1] @9
--
--tmp(30) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(31) := RET & "000" & "000000000"; -- RET
--
--tmp(32) := LDA & "001" & "000001000"; -- LDA [1] @8
--
--tmp(33) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(34) := CEQ & "010" & "000001110"; -- CEQ [2] @14
--
--tmp(35) := JEQ & "000" & "000100111"; -- JEQ @39
--
--tmp(36) := SOMA & "010" & "000001001"; -- SOMA [2] @9
--
--tmp(37) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(38) := RET & "000" & "000000000"; -- RET
--
--tmp(39) := LDA & "010" & "000001000"; -- LDA [2] @8
--
--tmp(40) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(41) := CEQ & "011" & "000001110"; -- CEQ [3] @14
--
--tmp(42) := JEQ & "000" & "000101110"; -- JEQ @46
--
--tmp(43) := SOMA & "011" & "000001001"; -- SOMA [3] @9
--
--tmp(44) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(45) := RET & "000" & "000000000"; -- RET
--
--tmp(46) := LDA & "011" & "000001000"; -- LDA [3] @8
--
--tmp(47) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(48) := CEQ & "100" & "000001110"; -- CEQ [4] @14
--
--tmp(49) := JEQ & "000" & "000110101"; -- JEQ @53
--
--tmp(50) := SOMA & "100" & "000001001"; -- SOMA [4] @9
--
--tmp(51) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(52) := RET & "000" & "000000000"; -- RET
--
--tmp(53) := LDA & "100" & "000001000"; -- LDA [4] @8
--
--tmp(54) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(55) := CEQ & "101" & "000001110"; -- CEQ [5] @14
--
--tmp(56) := JEQ & "000" & "000111100"; -- JEQ @60
--
--tmp(57) := SOMA & "101" & "000001001"; -- SOMA [5] @9
--
--tmp(58) := STA & "101" & "100100101"; -- STA [5] @293
--
--tmp(59) := RET & "000" & "000000000"; -- RET
--
--tmp(60) := LDI & "110" & "000000001"; -- LDI [6] $1
--
--tmp(61) := STA & "110" & "100000010"; -- STA [6] @258
--
--tmp(62) := RET & "000" & "000000000"; -- RET
--
--tmp(63) := LDI & "000" & "000000000"; -- LDI [0] $0
--
--tmp(64) := LDI & "001" & "000000000"; -- LDI [1] $0
--
--tmp(65) := LDI & "010" & "000000000"; -- LDI [2] $0
--
--tmp(66) := LDI & "011" & "000000000"; -- LDI [3] $0
--
--tmp(67) := LDI & "100" & "000000000"; -- LDI [4] $0
--
--tmp(68) := LDI & "101" & "000000000"; -- LDI [5] $0
--
--tmp(69) := STA & "000" & "100100000"; -- STA [0] @288
--
--tmp(70) := STA & "001" & "100100001"; -- STA [1] @289
--
--tmp(71) := STA & "010" & "100100010"; -- STA [2] @290
--
--tmp(72) := STA & "011" & "100100011"; -- STA [3] @291
--
--tmp(73) := STA & "100" & "100100100"; -- STA [4] @292
--
--tmp(74) := STA & "101" & "100100101"; -- STA [5] @293
--
--tmp(75) := JMP & "000" & "000001000"; -- JMP @8
--
--tmp(76) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(77) := STA & "110" & "100100000"; -- STA [6] @288
--
--tmp(78) := STA & "110" & "000000010"; -- STA [6] @2
--
--tmp(79) := STA & "000" & "111111110"; -- STA @510
--
--tmp(80) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(81) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(82) := JEQ & "000" & "001010000"; -- JEQ @80
--
--tmp(83) := STA & "000" & "111111110"; -- STA @510
--
--tmp(84) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(85) := STA & "110" & "100100001"; -- STA [6] @289
--
--tmp(86) := STA & "110" & "000000011"; -- STA [6] @3
--
--tmp(87) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(88) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(89) := JEQ & "000" & "001010111"; -- JEQ @87
--
--tmp(90) := STA & "000" & "111111110"; -- STA @510
--
--tmp(91) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(92) := STA & "110" & "100100010"; -- STA [6] @290
--
--tmp(93) := STA & "110" & "000000100"; -- STA [6] @4
--
--tmp(94) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(95) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(96) := JEQ & "000" & "001011110"; -- JEQ @94
--
--tmp(97) := STA & "000" & "111111110"; -- STA @510
--
--tmp(98) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(99) := STA & "110" & "100100011"; -- STA [6] @291
--
--tmp(100) := STA & "110" & "000000101"; -- STA [6] @5
--
--tmp(101) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(102) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(103) := JEQ & "000" & "001100101"; -- JEQ @101
--
--tmp(104) := STA & "000" & "111111110"; -- STA @510
--
--tmp(105) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(106) := STA & "110" & "100100100"; -- STA [6] @292
--
--tmp(107) := STA & "110" & "000000110"; -- STA [6] @6
--
--tmp(108) := LDA & "111" & "101100001"; -- LDA [7] @353
--
--tmp(109) := CEQ & "111" & "000001000"; -- CEQ [7] @8
--
--tmp(110) := JEQ & "000" & "001101100"; -- JEQ @108
--
--tmp(111) := STA & "000" & "111111110"; -- STA @510
--
--tmp(112) := LDA & "110" & "101000000"; -- LDA [6] @320
--
--tmp(113) := STA & "110" & "100100101"; -- STA [6] @293
--
--tmp(114) := STA & "110" & "000000111"; -- STA [6] @7
--
--tmp(115) := STA & "000" & "111111110"; -- STA @510
--
--tmp(116) := JMP & "000" & "000111111"; -- JMP @63



        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    data <= memROM (to_integer(unsigned(address)));
end architecture;