library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3;
			 opcodeSize: natural := 4
    );
   port (
          address : in std_logic_vector (addrWidth-1 DOWNTO 0);
          data : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;



architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDB : std_logic_vector(3 downto 0) := "1011";
  constant CLT  : std_logic_vector(3 downto 0) := "1100";
  constant JLT  : std_logic_vector(3 downto 0) := "1101";

  
  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin

tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(1) := STA & "111" & "000001000"; -- STA [7] @8

tmp(2) := LDI & "111" & "000000001"; -- LDI [7] $1

tmp(3) := STA & "111" & "000001001"; -- STA [7] @9

tmp(4) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(5) := STA & "111" & "000001011"; -- STA [7] @11

tmp(6) := LDI & "111" & "000001010"; -- LDI [7] $10

tmp(7) := STA & "111" & "000010010"; -- STA [7] @18

tmp(8) := LDI & "111" & "000001000"; -- LDI [7] $8

tmp(9) := STA & "111" & "000010110"; -- STA [7] @22

tmp(10) := LDI & "111" & "000001001"; -- LDI [7] $9

tmp(11) := STA & "111" & "000010001"; -- STA [7] @17

tmp(12) := STA & "111" & "000000010"; -- STA [7] @2

tmp(13) := STA & "111" & "000000100"; -- STA [7] @4

tmp(14) := STA & "111" & "000000110"; -- STA [7] @6

tmp(15) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(16) := STA & "111" & "000000111"; -- STA [7] @7

tmp(17) := LDI & "111" & "000000101"; -- LDI [7] $5

tmp(18) := STA & "111" & "000000011"; -- STA [7] @3

tmp(19) := STA & "111" & "000000101"; -- STA [7] @5

tmp(20) := LDI & "111" & "000000011"; -- LDI [7] $3

tmp(21) := STA & "111" & "000010011"; -- STA [7] @19

tmp(22) := STA & "000" & "111111111"; -- STA @511

tmp(23) := STA & "000" & "111111110"; -- STA @510

tmp(24) := JSR & "000" & "100101110"; -- JSR @302

tmp(25) := JMP & "000" & "010011101"; -- JMP @157

tmp(26) := LDA & "111" & "101100100"; -- LDA [7] @356

tmp(27) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(28) := JEQ & "000" & "010011101"; -- JEQ @157

tmp(29) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(30) := CEQ & "111" & "000001001"; -- CEQ [7] @9

tmp(31) := JEQ & "000" & "011011111"; -- JEQ @223

tmp(32) := LDA & "111" & "101100010"; -- LDA [7] @354

tmp(33) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(34) := JEQ & "000" & "001010001"; -- JEQ @81

tmp(35) := LDA & "111" & "101100011"; -- LDA [7] @355

tmp(36) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(37) := JEQ & "000" & "000101111"; -- JEQ @47

tmp(38) := LDA & "111" & "111111100"; -- LDA [7] @508

tmp(39) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(40) := STA & "000" & "111111101"; -- STA @509

tmp(41) := JEQ & "000" & "000011010"; -- JEQ @26

tmp(42) := JSR & "000" & "010111010"; -- JSR @186

tmp(43) := LDA & "110" & "000010100"; -- LDA [6] @20

tmp(44) := STA & "110" & "100000001"; -- STA [6] @257

tmp(45) := JSR & "000" & "001110000"; -- JSR @112

tmp(46) := JMP & "000" & "000011010"; -- JMP @26

tmp(47) := LDI & "110" & "000000000"; -- LDI [6] $0

tmp(48) := CEQ & "110" & "000010101"; -- CEQ [6] @21

tmp(49) := JEQ & "000" & "000111010"; -- JEQ @58

tmp(50) := LDI & "110" & "000000011"; -- LDI [6] $3

tmp(51) := STA & "110" & "000010011"; -- STA [6] @19

tmp(52) := LDI & "110" & "000000010"; -- LDI [6] $2

tmp(53) := STA & "110" & "000000111"; -- STA [6] @7

tmp(54) := LDA & "111" & "000010001"; -- LDA [7] @17

tmp(55) := STA & "111" & "000000110"; -- STA [7] @6

tmp(56) := JSR & "000" & "100101110"; -- JSR @302

tmp(57) := JSR & "000" & "000111101"; -- JSR @61

tmp(58) := JSR & "000" & "100110100"; -- JSR @308

tmp(59) := LDI & "111" & "000000100"; -- LDI [7] $4

tmp(60) := JMP & "000" & "100100010"; -- JMP @290

tmp(61) := LDA & "111" & "000010100"; -- LDA [7] @20

tmp(62) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(63) := JEQ & "000" & "100101011"; -- JEQ @299

tmp(64) := CEQ & "101" & "000001000"; -- CEQ [5] @8

tmp(65) := JEQ & "000" & "001000111"; -- JEQ @71

tmp(66) := LDI & "111" & "000000011"; -- LDI [7] $3

tmp(67) := STA & "111" & "000000110"; -- STA [7] @6

tmp(68) := SOMA & "100" & "000001011"; -- SOMA [4] @11

tmp(69) := SOMA & "101" & "000001001"; -- SOMA [5] @9

tmp(70) := RET & "000" & "000000000"; -- RET

tmp(71) := CLT & "100" & "000010110"; -- CLT [4] @22

tmp(72) := JLT & "000" & "001001110"; -- JLT @78

tmp(73) := LDI & "111" & "000000011"; -- LDI [7] $3

tmp(74) := STA & "111" & "000000110"; -- STA [7] @6

tmp(75) := LDA & "101" & "000001011"; -- LDA [5] @11

tmp(76) := SUB & "100" & "000010110"; -- SUB [4] @22

tmp(77) := RET & "000" & "000000000"; -- RET

tmp(78) := SOMA & "100" & "000001011"; -- SOMA [4] @11

tmp(79) := LDA & "101" & "000001001"; -- LDA [5] @9

tmp(80) := RET & "000" & "000000000"; -- RET

tmp(81) := LDI & "110" & "000000001"; -- LDI [6] $1

tmp(82) := CEQ & "110" & "000010101"; -- CEQ [6] @21

tmp(83) := JEQ & "000" & "001011000"; -- JEQ @88

tmp(84) := STA & "110" & "000010011"; -- STA [6] @19

tmp(85) := STA & "110" & "000000111"; -- STA [6] @7

tmp(86) := JSR & "000" & "001011010"; -- JSR @90

tmp(87) := JSR & "000" & "100110001"; -- JSR @305

tmp(88) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(89) := JMP & "000" & "100100010"; -- JMP @290

tmp(90) := CEQ & "101" & "000001000"; -- CEQ [5] @8

tmp(91) := JEQ & "000" & "100101011"; -- JEQ @299

tmp(92) := CEQ & "101" & "000001001"; -- CEQ [5] @9

tmp(93) := JEQ & "000" & "001100101"; -- JEQ @101

tmp(94) := CLT & "100" & "000001011"; -- CLT [4] @11

tmp(95) := JLT & "000" & "001101010"; -- JLT @106

tmp(96) := SUB & "101" & "000001001"; -- SUB [5] @9

tmp(97) := SUB & "100" & "000001011"; -- SUB [4] @11

tmp(98) := LDA & "111" & "000001001"; -- LDA [7] @9

tmp(99) := STA & "111" & "000000110"; -- STA [7] @6

tmp(100) := JMP & "000" & "100110111"; -- JMP @311

tmp(101) := CLT & "100" & "000001011"; -- CLT [4] @11

tmp(102) := JLT & "000" & "100101011"; -- JLT @299

tmp(103) := SUB & "100" & "000001011"; -- SUB [4] @11

tmp(104) := LDA & "101" & "000001000"; -- LDA [5] @8

tmp(105) := JMP & "000" & "100110111"; -- JMP @311

tmp(106) := SUB & "100" & "000001011"; -- SUB [4] @11

tmp(107) := SOMA & "100" & "000010010"; -- SOMA [4] @18

tmp(108) := LDA & "101" & "000001000"; -- LDA [5] @8

tmp(109) := LDA & "111" & "000010001"; -- LDA [7] @17

tmp(110) := STA & "111" & "000000110"; -- STA [7] @6

tmp(111) := JMP & "000" & "100110111"; -- JMP @311

tmp(112) := CEQ & "000" & "000000010"; -- CEQ [0] @2

tmp(113) := JEQ & "000" & "001110101"; -- JEQ @117

tmp(114) := SOMA & "000" & "000001001"; -- SOMA [0] @9

tmp(115) := STA & "000" & "100100000"; -- STA [0] @288

tmp(116) := RET & "000" & "000000000"; -- RET

tmp(117) := LDA & "000" & "000001000"; -- LDA [0] @8

tmp(118) := STA & "000" & "100100000"; -- STA [0] @288

tmp(119) := CEQ & "001" & "000000011"; -- CEQ [1] @3

tmp(120) := JEQ & "000" & "001111100"; -- JEQ @124

tmp(121) := SOMA & "001" & "000001001"; -- SOMA [1] @9

tmp(122) := STA & "001" & "100100001"; -- STA [1] @289

tmp(123) := RET & "000" & "000000000"; -- RET

tmp(124) := LDA & "001" & "000001000"; -- LDA [1] @8

tmp(125) := STA & "001" & "100100001"; -- STA [1] @289

tmp(126) := CEQ & "010" & "000000100"; -- CEQ [2] @4

tmp(127) := JEQ & "000" & "010000011"; -- JEQ @131

tmp(128) := SOMA & "010" & "000001001"; -- SOMA [2] @9

tmp(129) := STA & "010" & "100100010"; -- STA [2] @290

tmp(130) := RET & "000" & "000000000"; -- RET

tmp(131) := LDA & "010" & "000001000"; -- LDA [2] @8

tmp(132) := STA & "010" & "100100010"; -- STA [2] @290

tmp(133) := CEQ & "011" & "000000101"; -- CEQ [3] @5

tmp(134) := JEQ & "000" & "010001010"; -- JEQ @138

tmp(135) := SOMA & "011" & "000001001"; -- SOMA [3] @9

tmp(136) := STA & "011" & "100100011"; -- STA [3] @291

tmp(137) := RET & "000" & "000000000"; -- RET

tmp(138) := LDA & "011" & "000001000"; -- LDA [3] @8

tmp(139) := STA & "011" & "100100011"; -- STA [3] @291

tmp(140) := CEQ & "100" & "000000110"; -- CEQ [4] @6

tmp(141) := JEQ & "000" & "010010001"; -- JEQ @145

tmp(142) := SOMA & "100" & "000001001"; -- SOMA [4] @9

tmp(143) := STA & "100" & "100100100"; -- STA [4] @292

tmp(144) := RET & "000" & "000000000"; -- RET

tmp(145) := LDA & "100" & "000001000"; -- LDA [4] @8

tmp(146) := STA & "100" & "100100100"; -- STA [4] @292

tmp(147) := CEQ & "101" & "000000111"; -- CEQ [5] @7

tmp(148) := JEQ & "000" & "010100111"; -- JEQ @167

tmp(149) := SOMA & "101" & "000001001"; -- SOMA [5] @9

tmp(150) := STA & "101" & "100100101"; -- STA [5] @293

tmp(151) := CEQ & "101" & "000000111"; -- CEQ [5] @7

tmp(152) := JEQ & "000" & "010011010"; -- JEQ @154

tmp(153) := RET & "000" & "000000000"; -- RET

tmp(154) := LDA & "111" & "000010011"; -- LDA [7] @19

tmp(155) := STA & "111" & "000000110"; -- STA [7] @6

tmp(156) := RET & "000" & "000000000"; -- RET

tmp(157) := LDI & "111" & "000001001"; -- LDI [7] $9

tmp(158) := STA & "111" & "000000110"; -- STA [7] @6

tmp(159) := LDI & "000" & "000000000"; -- LDI [0] $0

tmp(160) := LDI & "001" & "000000000"; -- LDI [1] $0

tmp(161) := LDI & "010" & "000000000"; -- LDI [2] $0

tmp(162) := LDI & "011" & "000000000"; -- LDI [3] $0

tmp(163) := LDI & "100" & "000000000"; -- LDI [4] $0

tmp(164) := LDI & "101" & "000000000"; -- LDI [5] $0

tmp(165) := JSR & "000" & "010111010"; -- JSR @186

tmp(166) := JMP & "000" & "000011010"; -- JMP @26

tmp(167) := LDI & "111" & "000001001"; -- LDI [7] $9

tmp(168) := STA & "111" & "000000110"; -- STA [7] @6

tmp(169) := LDI & "000" & "000000000"; -- LDI [0] $0

tmp(170) := LDI & "001" & "000000000"; -- LDI [1] $0

tmp(171) := LDI & "010" & "000000000"; -- LDI [2] $0

tmp(172) := LDI & "011" & "000000000"; -- LDI [3] $0

tmp(173) := LDI & "100" & "000000000"; -- LDI [4] $0

tmp(174) := STA & "101" & "000001101"; -- STA [5] @13

tmp(175) := LDA & "110" & "000001101"; -- LDA [6] @13

tmp(176) := LDI & "101" & "000000000"; -- LDI [5] $0

tmp(177) := JSR & "000" & "010111010"; -- JSR @186

tmp(178) := CEQ & "110" & "000001011"; -- CEQ [6] @11

tmp(179) := JEQ & "000" & "000011010"; -- JEQ @26

tmp(180) := JSR & "000" & "010110110"; -- JSR @182

tmp(181) := JMP & "000" & "000011010"; -- JMP @26

tmp(182) := LDA & "111" & "000010100"; -- LDA [7] @20

tmp(183) := SOMA & "111" & "000001001"; -- SOMA [7] @9

tmp(184) := ANDB & "111" & "000001001"; -- ANDB [7] @9

tmp(185) := STA & "111" & "000010100"; -- STA [7] @20

tmp(186) := STA & "000" & "100100000"; -- STA [0] @288

tmp(187) := STA & "001" & "100100001"; -- STA [1] @289

tmp(188) := STA & "010" & "100100010"; -- STA [2] @290

tmp(189) := STA & "011" & "100100011"; -- STA [3] @291

tmp(190) := STA & "100" & "100100100"; -- STA [4] @292

tmp(191) := STA & "101" & "100100101"; -- STA [5] @293

tmp(192) := RET & "000" & "000000000"; -- RET

tmp(193) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(194) := STA & "111" & "100100000"; -- STA [7] @288

tmp(195) := STA & "111" & "100100001"; -- STA [7] @289

tmp(196) := STA & "111" & "100100010"; -- STA [7] @290

tmp(197) := STA & "111" & "100100011"; -- STA [7] @291

tmp(198) := STA & "111" & "100100100"; -- STA [7] @292

tmp(199) := STA & "111" & "100100101"; -- STA [7] @293

tmp(200) := RET & "000" & "000000000"; -- RET

tmp(201) := JSR & "000" & "011000001"; -- JSR @193

tmp(202) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(203) := LDA & "111" & "000000010"; -- LDA [7] @2

tmp(204) := JSR & "000" & "100011010"; -- JSR @282

tmp(205) := STA & "110" & "100100000"; -- STA [6] @288

tmp(206) := STA & "110" & "000001100"; -- STA [6] @12

tmp(207) := LDA & "000" & "000001100"; -- LDA [0] @12

tmp(208) := STA & "000" & "111111110"; -- STA @510

tmp(209) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(210) := STA & "111" & "100000000"; -- STA [7] @256

tmp(211) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(212) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(213) := JEQ & "000" & "011010011"; -- JEQ @211

tmp(214) := STA & "000" & "111111110"; -- STA @510

tmp(215) := LDI & "111" & "000000100"; -- LDI [7] $4

tmp(216) := STA & "111" & "100000000"; -- STA [7] @256

tmp(217) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(218) := LDA & "111" & "000000011"; -- LDA [7] @3

tmp(219) := JSR & "000" & "100011010"; -- JSR @282

tmp(220) := STA & "110" & "100100001"; -- STA [6] @289

tmp(221) := STA & "110" & "000001100"; -- STA [6] @12

tmp(222) := LDA & "001" & "000001100"; -- LDA [1] @12

tmp(223) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(224) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(225) := JEQ & "000" & "011011111"; -- JEQ @223

tmp(226) := STA & "000" & "111111110"; -- STA @510

tmp(227) := LDI & "111" & "000001000"; -- LDI [7] $8

tmp(228) := STA & "111" & "100000000"; -- STA [7] @256

tmp(229) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(230) := LDA & "111" & "000000100"; -- LDA [7] @4

tmp(231) := JSR & "000" & "100011010"; -- JSR @282

tmp(232) := STA & "110" & "100100010"; -- STA [6] @290

tmp(233) := STA & "110" & "000001100"; -- STA [6] @12

tmp(234) := LDA & "010" & "000001100"; -- LDA [2] @12

tmp(235) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(236) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(237) := JEQ & "000" & "011101011"; -- JEQ @235

tmp(238) := STA & "000" & "111111110"; -- STA @510

tmp(239) := LDI & "111" & "000010000"; -- LDI [7] $16

tmp(240) := STA & "111" & "100000000"; -- STA [7] @256

tmp(241) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(242) := LDA & "111" & "000000101"; -- LDA [7] @5

tmp(243) := JSR & "000" & "100011010"; -- JSR @282

tmp(244) := STA & "110" & "100100011"; -- STA [6] @291

tmp(245) := STA & "110" & "000001100"; -- STA [6] @12

tmp(246) := LDA & "011" & "000001100"; -- LDA [3] @12

tmp(247) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(248) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(249) := JEQ & "000" & "011110111"; -- JEQ @247

tmp(250) := STA & "000" & "111111110"; -- STA @510

tmp(251) := LDI & "111" & "000100000"; -- LDI [7] $32

tmp(252) := STA & "111" & "100000000"; -- STA [7] @256

tmp(253) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(254) := LDA & "111" & "000000110"; -- LDA [7] @6

tmp(255) := JSR & "000" & "100011010"; -- JSR @282

tmp(256) := STA & "110" & "100100100"; -- STA [6] @292

tmp(257) := STA & "110" & "000001100"; -- STA [6] @12

tmp(258) := LDA & "100" & "000001100"; -- LDA [4] @12

tmp(259) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(260) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(261) := JEQ & "000" & "100000011"; -- JEQ @259

tmp(262) := STA & "000" & "111111110"; -- STA @510

tmp(263) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(264) := STA & "111" & "100000000"; -- STA [7] @256

tmp(265) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(266) := LDA & "111" & "000000111"; -- LDA [7] @7

tmp(267) := JSR & "000" & "100011010"; -- JSR @282

tmp(268) := STA & "110" & "100100101"; -- STA [6] @293

tmp(269) := STA & "110" & "000001100"; -- STA [6] @12

tmp(270) := LDA & "101" & "000001100"; -- LDA [5] @12

tmp(271) := CLT & "110" & "000000111"; -- CLT [6] @7

tmp(272) := JLT & "000" & "100010100"; -- JLT @276

tmp(273) := LDA & "100" & "000010011"; -- LDA [4] @19

tmp(274) := STA & "100" & "100100100"; -- STA [4] @292

tmp(275) := STA & "100" & "000000110"; -- STA [4] @6

tmp(276) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(277) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(278) := JEQ & "000" & "100010100"; -- JEQ @276

tmp(279) := STA & "000" & "111111110"; -- STA @510

tmp(280) := JSR & "000" & "010111010"; -- JSR @186

tmp(281) := JMP & "000" & "000011010"; -- JMP @26

tmp(282) := STA & "111" & "000001101"; -- STA [7] @13

tmp(283) := CLT & "110" & "000001101"; -- CLT [6] @13

tmp(284) := JLT & "000" & "100100000"; -- JLT @288

tmp(285) := LDA & "110" & "000001101"; -- LDA [6] @13

tmp(286) := LDA & "111" & "000001001"; -- LDA [7] @9

tmp(287) := RET & "000" & "000000000"; -- RET

tmp(288) := LDA & "111" & "000001000"; -- LDA [7] @8

tmp(289) := RET & "000" & "000000000"; -- RET

tmp(290) := LDA & "110" & "000001000"; -- LDA [6] @8

tmp(291) := STA & "110" & "100100000"; -- STA [6] @288

tmp(292) := STA & "110" & "100100001"; -- STA [6] @289

tmp(293) := STA & "110" & "100100010"; -- STA [6] @290

tmp(294) := STA & "110" & "100100011"; -- STA [6] @291

tmp(295) := STA & "111" & "100100100"; -- STA [7] @292

tmp(296) := LDA & "111" & "000000111"; -- LDA [7] @7

tmp(297) := STA & "111" & "100100101"; -- STA [7] @293

tmp(298) := JMP & "000" & "000011010"; -- JMP @26

tmp(299) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(300) := STA & "111" & "000010100"; -- STA [7] @20

tmp(301) := RET & "000" & "000000000"; -- RET

tmp(302) := LDA & "110" & "000001000"; -- LDA [6] @8

tmp(303) := STA & "110" & "000010101"; -- STA [6] @21

tmp(304) := RET & "000" & "000000000"; -- RET

tmp(305) := LDA & "110" & "000001001"; -- LDA [6] @9

tmp(306) := STA & "110" & "000010101"; -- STA [6] @21

tmp(307) := RET & "000" & "000000000"; -- RET

tmp(308) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(309) := STA & "111" & "000010100"; -- STA [7] @20

tmp(310) := RET & "000" & "000000000"; -- RET

tmp(311) := LDI & "111" & "000000001"; -- LDI [7] $1

tmp(312) := STA & "111" & "000010100"; -- STA [7] @20

tmp(313) := RET & "000" & "000000000"; -- RET

        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    data <= memROM (to_integer(unsigned(address)));
end architecture;