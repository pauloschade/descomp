library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 3;
			 opcodeSize: natural := 4
    );
   port (
          address : in std_logic_vector (addrWidth-1 DOWNTO 0);
          data : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;



architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDB : std_logic_vector(3 downto 0) := "1011";
  constant CLT  : std_logic_vector(3 downto 0) := "1100";
  constant JLT  : std_logic_vector(3 downto 0) := "1101";

  
  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin

 tmp(0) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(1) := STA & "111" & "000001000"; -- STA [7] @8

tmp(2) := LDI & "111" & "000000001"; -- LDI [7] $1

tmp(3) := STA & "111" & "000001001"; -- STA [7] @9

tmp(4) := LDI & "111" & "000001001"; -- LDI [7] $9

tmp(5) := STA & "111" & "000010001"; -- STA [7] @17

tmp(6) := STA & "111" & "000000010"; -- STA [7] @2

tmp(7) := STA & "111" & "000000100"; -- STA [7] @4

tmp(8) := STA & "111" & "000000110"; -- STA [7] @6

tmp(9) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(10) := STA & "111" & "000000111"; -- STA [7] @7

tmp(11) := LDI & "111" & "000000101"; -- LDI [7] $5

tmp(12) := STA & "111" & "000000011"; -- STA [7] @3

tmp(13) := STA & "111" & "000000101"; -- STA [7] @5

tmp(14) := LDI & "111" & "000000011"; -- LDI [7] $3

tmp(15) := STA & "111" & "000010010"; -- STA [7] @18

tmp(16) := STA & "000" & "111111111"; -- STA @511

tmp(17) := STA & "000" & "111111110"; -- STA @510

tmp(18) := JMP & "000" & "001100001"; -- JMP @97

tmp(19) := LDA & "111" & "101100100"; -- LDA [7] @356

tmp(20) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(21) := JEQ & "000" & "001100001"; -- JEQ @97

tmp(22) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(23) := CEQ & "111" & "000001001"; -- CEQ [7] @9

tmp(24) := JEQ & "000" & "010010000"; -- JEQ @144

tmp(25) := LDA & "111" & "101100010"; -- LDA [7] @354

tmp(26) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(27) := JEQ & "000" & "000101110"; -- JEQ @46

tmp(28) := LDA & "111" & "101100011"; -- LDA [7] @355

tmp(29) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(30) := JEQ & "000" & "000101000"; -- JEQ @40

tmp(31) := LDA & "111" & "101100000"; -- LDA [7] @352

tmp(32) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(33) := JEQ & "000" & "000010011"; -- JEQ @19

tmp(34) := JSR & "000" & "001101011"; -- JSR @107

tmp(35) := LDA & "110" & "000001000"; -- LDA [6] @8

tmp(36) := STA & "110" & "100000001"; -- STA [6] @257

tmp(37) := STA & "000" & "111111111"; -- STA @511

tmp(38) := JSR & "000" & "001000111"; -- JSR @71

tmp(39) := JMP & "000" & "000010011"; -- JMP @19

tmp(40) := LDI & "110" & "000000011"; -- LDI [6] $3

tmp(41) := STA & "110" & "000010010"; -- STA [6] @18

tmp(42) := LDI & "110" & "000000010"; -- LDI [6] $2

tmp(43) := STA & "110" & "000000111"; -- STA [6] @7

tmp(44) := LDI & "111" & "000000100"; -- LDI [7] $4

tmp(45) := JMP & "000" & "011001110"; -- JMP @206

tmp(46) := LDI & "110" & "000000001"; -- LDI [6] $1

tmp(47) := STA & "110" & "000010010"; -- STA [6] @18

tmp(48) := LDI & "110" & "000000001"; -- LDI [6] $1

tmp(49) := STA & "110" & "000000111"; -- STA [6] @7

tmp(50) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(51) := JMP & "000" & "011001110"; -- JMP @206

tmp(52) := CEQ & "000" & "000000010"; -- CEQ [0] @2

tmp(53) := JEQ & "000" & "000111001"; -- JEQ @57

tmp(54) := SOMA & "000" & "000001001"; -- SOMA [0] @9

tmp(55) := STA & "000" & "100100000"; -- STA [0] @288

tmp(56) := RET & "000" & "000000000"; -- RET

tmp(57) := LDA & "000" & "000001000"; -- LDA [0] @8

tmp(58) := STA & "000" & "100100000"; -- STA [0] @288

tmp(59) := CEQ & "001" & "000000011"; -- CEQ [1] @3

tmp(60) := JEQ & "000" & "001000000"; -- JEQ @64

tmp(61) := SOMA & "001" & "000001001"; -- SOMA [1] @9

tmp(62) := STA & "001" & "100100001"; -- STA [1] @289

tmp(63) := RET & "000" & "000000000"; -- RET

tmp(64) := LDA & "001" & "000001000"; -- LDA [1] @8

tmp(65) := STA & "001" & "100100001"; -- STA [1] @289

tmp(66) := CEQ & "010" & "000000100"; -- CEQ [2] @4

tmp(67) := JEQ & "000" & "001000111"; -- JEQ @71

tmp(68) := SOMA & "010" & "000001001"; -- SOMA [2] @9

tmp(69) := STA & "010" & "100100010"; -- STA [2] @290

tmp(70) := RET & "000" & "000000000"; -- RET

tmp(71) := LDA & "010" & "000001000"; -- LDA [2] @8

tmp(72) := STA & "010" & "100100010"; -- STA [2] @290

tmp(73) := CEQ & "011" & "000000101"; -- CEQ [3] @5

tmp(74) := JEQ & "000" & "001001110"; -- JEQ @78

tmp(75) := SOMA & "011" & "000001001"; -- SOMA [3] @9

tmp(76) := STA & "011" & "100100011"; -- STA [3] @291

tmp(77) := RET & "000" & "000000000"; -- RET

tmp(78) := LDA & "011" & "000001000"; -- LDA [3] @8

tmp(79) := STA & "011" & "100100011"; -- STA [3] @291

tmp(80) := CEQ & "100" & "000000110"; -- CEQ [4] @6

tmp(81) := JEQ & "000" & "001010101"; -- JEQ @85

tmp(82) := SOMA & "100" & "000001001"; -- SOMA [4] @9

tmp(83) := STA & "100" & "100100100"; -- STA [4] @292

tmp(84) := RET & "000" & "000000000"; -- RET

tmp(85) := LDA & "100" & "000001000"; -- LDA [4] @8

tmp(86) := STA & "100" & "100100100"; -- STA [4] @292

tmp(87) := CEQ & "101" & "000000111"; -- CEQ [5] @7

tmp(88) := JEQ & "000" & "001100001"; -- JEQ @97

tmp(89) := SOMA & "101" & "000001001"; -- SOMA [5] @9

tmp(90) := STA & "101" & "100100101"; -- STA [5] @293

tmp(91) := CEQ & "101" & "000000111"; -- CEQ [5] @7

tmp(92) := JEQ & "000" & "001011110"; -- JEQ @94

tmp(93) := RET & "000" & "000000000"; -- RET

tmp(94) := LDA & "111" & "000010010"; -- LDA [7] @18

tmp(95) := STA & "111" & "000000110"; -- STA [7] @6

tmp(96) := RET & "000" & "000000000"; -- RET

tmp(97) := LDI & "111" & "000001001"; -- LDI [7] $9

tmp(98) := STA & "111" & "000000110"; -- STA [7] @6

tmp(99) := LDI & "000" & "000000000"; -- LDI [0] $0

tmp(100) := LDI & "001" & "000000000"; -- LDI [1] $0

tmp(101) := LDI & "010" & "000000000"; -- LDI [2] $0

tmp(102) := LDI & "011" & "000000000"; -- LDI [3] $0

tmp(103) := LDI & "100" & "000000000"; -- LDI [4] $0

tmp(104) := LDI & "101" & "000000000"; -- LDI [5] $0

tmp(105) := JSR & "000" & "001101011"; -- JSR @107

tmp(106) := JMP & "000" & "000010011"; -- JMP @19

tmp(107) := STA & "000" & "100100000"; -- STA [0] @288

tmp(108) := STA & "001" & "100100001"; -- STA [1] @289

tmp(109) := STA & "010" & "100100010"; -- STA [2] @290

tmp(110) := STA & "011" & "100100011"; -- STA [3] @291

tmp(111) := STA & "100" & "100100100"; -- STA [4] @292

tmp(112) := STA & "101" & "100100101"; -- STA [5] @293

tmp(113) := RET & "000" & "000000000"; -- RET

tmp(114) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(115) := STA & "111" & "100100000"; -- STA [7] @288

tmp(116) := STA & "111" & "100100001"; -- STA [7] @289

tmp(117) := STA & "111" & "100100010"; -- STA [7] @290

tmp(118) := STA & "111" & "100100011"; -- STA [7] @291

tmp(119) := STA & "111" & "100100100"; -- STA [7] @292

tmp(120) := STA & "111" & "100100101"; -- STA [7] @293

tmp(121) := RET & "000" & "000000000"; -- RET

tmp(122) := JSR & "000" & "001110010"; -- JSR @114

tmp(123) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(124) := LDA & "111" & "000000010"; -- LDA [7] @2

tmp(125) := JSR & "000" & "011000110"; -- JSR @198

tmp(126) := STA & "110" & "100100000"; -- STA [6] @288

tmp(127) := STA & "110" & "000001100"; -- STA [6] @12

tmp(128) := LDA & "000" & "000001100"; -- LDA [0] @12

tmp(129) := STA & "000" & "111111110"; -- STA @510

tmp(130) := LDI & "111" & "000000010"; -- LDI [7] $2

tmp(131) := STA & "111" & "100000000"; -- STA [7] @256

tmp(132) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(133) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(134) := JEQ & "000" & "010000100"; -- JEQ @132

tmp(135) := STA & "000" & "111111110"; -- STA @510

tmp(136) := LDI & "111" & "000000100"; -- LDI [7] $4

tmp(137) := STA & "111" & "100000000"; -- STA [7] @256

tmp(138) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(139) := LDA & "111" & "000000011"; -- LDA [7] @3

tmp(140) := JSR & "000" & "011000110"; -- JSR @198

tmp(141) := STA & "110" & "100100001"; -- STA [6] @289

tmp(142) := STA & "110" & "000001100"; -- STA [6] @12

tmp(143) := LDA & "001" & "000001100"; -- LDA [1] @12

tmp(144) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(145) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(146) := JEQ & "000" & "010010000"; -- JEQ @144

tmp(147) := STA & "000" & "111111110"; -- STA @510

tmp(148) := LDI & "111" & "000001000"; -- LDI [7] $8

tmp(149) := STA & "111" & "100000000"; -- STA [7] @256

tmp(150) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(151) := LDA & "111" & "000000100"; -- LDA [7] @4

tmp(152) := JSR & "000" & "011000110"; -- JSR @198

tmp(153) := STA & "110" & "100100010"; -- STA [6] @290

tmp(154) := STA & "110" & "000001100"; -- STA [6] @12

tmp(155) := LDA & "010" & "000001100"; -- LDA [2] @12

tmp(156) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(157) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(158) := JEQ & "000" & "010011100"; -- JEQ @156

tmp(159) := STA & "000" & "111111110"; -- STA @510

tmp(160) := LDI & "111" & "000010000"; -- LDI [7] $16

tmp(161) := STA & "111" & "100000000"; -- STA [7] @256

tmp(162) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(163) := LDA & "111" & "000000101"; -- LDA [7] @5

tmp(164) := JSR & "000" & "011000110"; -- JSR @198

tmp(165) := STA & "110" & "100100011"; -- STA [6] @291

tmp(166) := STA & "110" & "000001100"; -- STA [6] @12

tmp(167) := LDA & "011" & "000001100"; -- LDA [3] @12

tmp(168) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(169) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(170) := JEQ & "000" & "010101000"; -- JEQ @168

tmp(171) := STA & "000" & "111111110"; -- STA @510

tmp(172) := LDI & "111" & "000100000"; -- LDI [7] $32

tmp(173) := STA & "111" & "100000000"; -- STA [7] @256

tmp(174) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(175) := LDA & "111" & "000000110"; -- LDA [7] @6

tmp(176) := JSR & "000" & "011000110"; -- JSR @198

tmp(177) := STA & "110" & "100100100"; -- STA [6] @292

tmp(178) := STA & "110" & "000001100"; -- STA [6] @12

tmp(179) := LDA & "100" & "000001100"; -- LDA [4] @12

tmp(180) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(181) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(182) := JEQ & "000" & "010110100"; -- JEQ @180

tmp(183) := STA & "000" & "111111110"; -- STA @510

tmp(184) := LDI & "111" & "000000000"; -- LDI [7] $0

tmp(185) := STA & "111" & "100000000"; -- STA [7] @256

tmp(186) := LDA & "110" & "101000000"; -- LDA [6] @320

tmp(187) := LDA & "111" & "000000111"; -- LDA [7] @7

tmp(188) := JSR & "000" & "011000110"; -- JSR @198

tmp(189) := STA & "110" & "100100101"; -- STA [6] @293

tmp(190) := STA & "110" & "000001100"; -- STA [6] @12

tmp(191) := LDA & "101" & "000001100"; -- LDA [5] @12

tmp(192) := LDA & "111" & "101100001"; -- LDA [7] @353

tmp(193) := CEQ & "111" & "000001000"; -- CEQ [7] @8

tmp(194) := JEQ & "000" & "011000000"; -- JEQ @192

tmp(195) := STA & "000" & "111111110"; -- STA @510

tmp(196) := JSR & "000" & "001101011"; -- JSR @107

tmp(197) := JMP & "000" & "000010011"; -- JMP @19

tmp(198) := STA & "111" & "000001101"; -- STA [7] @13

tmp(199) := CLT & "110" & "000001101"; -- CLT [6] @13

tmp(200) := JLT & "000" & "011001100"; -- JLT @204

tmp(201) := LDA & "110" & "000001101"; -- LDA [6] @13

tmp(202) := LDA & "111" & "000001001"; -- LDA [7] @9

tmp(203) := RET & "000" & "000000000"; -- RET

tmp(204) := LDA & "111" & "000001000"; -- LDA [7] @8

tmp(205) := RET & "000" & "000000000"; -- RET

tmp(206) := LDA & "110" & "000001000"; -- LDA [6] @8

tmp(207) := STA & "110" & "100100000"; -- STA [6] @288

tmp(208) := STA & "110" & "100100001"; -- STA [6] @289

tmp(209) := STA & "110" & "100100010"; -- STA [6] @290

tmp(210) := STA & "110" & "100100011"; -- STA [6] @291

tmp(211) := STA & "111" & "100100100"; -- STA [7] @292

tmp(212) := LDA & "111" & "000000111"; -- LDA [7] @7

tmp(213) := STA & "111" & "100100101"; -- STA [7] @293

tmp(214) := JMP & "000" & "000010011"; -- JMP @19

  
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    data <= memROM (to_integer(unsigned(address)));
end architecture;